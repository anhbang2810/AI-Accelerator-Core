// =============================================================================
// Module:      tb_npu_pe (Unit Test)
// Description: Kiem thu (ALU) nap tay
// =============================================================================
`timescale 1ns/1ps

module tb_npu_pe;

  parameter DATA_WIDTH = 8;
  parameter ACC_WIDTH  = 20;

  logic clk = 0;
  logic rst_n = 0;
  
  logic i_valid = 0;
  logic i_last = 0;
  logic signed [DATA_WIDTH-1:0] i_feature;
  logic signed [DATA_WIDTH-1:0] i_weight;
  logic signed [ACC_WIDTH-1:0]  i_bias;
  
  logic o_valid;
  logic signed [DATA_WIDTH-1:0] o_result;

  npu_pe #(
    .DATA_WIDTH(DATA_WIDTH),
    .ACC_WIDTH(ACC_WIDTH)
  ) DUT (
    .clk(clk),
    .rst_n(rst_n),
    .i_valid(i_valid),
    .i_last(i_last),
    .i_feature(i_feature),
    .i_weight(i_weight),
    .i_bias(i_bias),
    .o_valid(o_valid),
    .o_result(o_result)
  );

  always #5 clk = ~clk;

  // ---------------------------------------------------------------------------
  // TASK: Gui goi du lieu (Helper Function)
  // ---------------------------------------------------------------------------
  task send_packet(
    input signed [DATA_WIDTH-1:0] feat, 
    input signed [DATA_WIDTH-1:0] w, 
    input is_end
  );
    begin
      @(posedge clk); 
      i_valid   <= 1;
      i_feature <= feat;
      i_weight  <= w;
      i_last    <= is_end;
    end
  endtask

  initial begin
    $display("==================================================");
    $display("   STARTING UNIT TEST: NPU PROCESSING ELEMENT     ");
    $display("==================================================");

    // --- B1 - Reset ---
    rst_n = 0; i_bias = 0;
    #20 rst_n = 1;

    // --- TEST CASE 1: Tinh toan so Duong (Normal Operation) ---
    // ReLU( (10*2) + (5*-3) + (2*4) + 5 ) = 18
    $display("\n[TEST 1] Testing MAC operation (Positive Output)...");
    
    i_bias = 5; 
    // Burst
    send_packet(8'd10,  8'd2,  0); // 10 * 2
    send_packet(8'd5,  -8'd3,  0); // 5 * -3
    send_packet(8'd2,   8'd4,  1); // 2 * 4 (i_last = 1)

    // Ngat tin hieu sau khi gui xong
    @(posedge clk);
    i_valid <= 0; i_last <= 0; i_feature <= 0; i_weight <= 0;

    // Cho ket qua
    wait(o_valid);
    @(negedge clk); 

    if (o_result === 8'd18) 
      $display(">> RESULT: %d (Expected: 18) -> PASS [OK]", o_result);
    else 
      $display(">> RESULT: %d (Expected: 18) -> FAIL [X]", o_result);

    
    // --- TEST CASE 2: Tinh so am (ReLU Check) ---
    // ReLU( (2*-10) + 5 ) = ReLU(-15) = 0
    #30; 
    $display("\n[TEST 2] Testing ReLU Activation (Negative Input)...");
    
    i_bias = 5;
    send_packet(8'd2, -8'd10, 1); // Gui 1 goi du lieu

    @(posedge clk);
    i_valid <= 0; i_last <= 0;

    wait(o_valid);
    @(negedge clk);

    if (o_result === 8'd0) 
      $display(">> RESULT: %d (Expected: 0 - ReLU Active) -> PASS [OK]", o_result);
    else 
      $display(">> RESULT: %d (Expected: 0) -> FAIL [X]", o_result);

    #50;
    $display("==================================================");
    $display("   UNIT TEST FINISHED                             ");
    $display("==================================================");
    $stop;
  end

endmodule